module parity_generator(



);


endmodule